-- author: R.D. Beyers
-- updated on 29/04/2015
-- STELLENBOSCH UNIVERSITY

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY CLK_SOURCE IS
	PORT
	(
		CLOCK_50	:	IN STD_LOGIC; -- the 50 MHz clock source on the DE0 board
		CPU_CLK		:	OUT STD_LOGIC -- the cpu clock source
	);
END CLK_SOURCE;

ARCHITECTURE STRUCTURE OF CLK_SOURCE IS	
	SIGNAL CPU_CLK_SIG	:	STD_LOGIC;
BEGIN
	CPU_CLK <= CPU_CLK_SIG;	
	PROCESS (CLOCK_50)
		VARIABLE CPU_CLK_CNT  : INTEGER RANGE 0 TO 50000000;
	BEGIN
		-- Generate CPU clock by dividing the 50 MHz clock by 2*CPU_CLK_CNT
		IF CLOCK_50'EVENT AND CLOCK_50 = '1' THEN
			CPU_CLK_CNT := CPU_CLK_CNT + 1;
			IF CPU_CLK_CNT = 25000000 THEN
				CPU_CLK_CNT := 0;
				CPU_CLK_SIG <= NOT CPU_CLK_SIG;
			END IF;
		END IF;
	END PROCESS;
END STRUCTURE;
